LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY PWM1 IS 
PORT(
		ENTRADA_RELOJ: IN STD_LOGIC;
		SELECTOR: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		SALIDA_PWM: OUT STD_LOGIC
	 );
END PWM1;

ARCHITECTURE MODULACION OF PWM1 IS 
SIGNAL CUENTA: STD_LOGIC_VECTOR (3 DOWNTO 0):= "0000";
BEGIN
   PROCESS (ENTRADA_RELOJ) 
	BEGIN 
		IF (ENTRADA_RELOJ'EVENT AND ENTRADA_RELOJ = '0') THEN --Preguntamos por la entrada de reloj y si está en 1 
		CUENTA <= CUENTA + "0001";
		END IF;
	END PROCESS;
	
	WITH SELECTOR SELECT  --USAMOS EL SELECTOR PARA MOSTRAR EL BIT DETERMINADO DE UNA CUENTA 
	
	SALIDA_PWM <= CUENTA(0) WHEN "00", --ELEGIMOS QUE LA SALIDA DEL PWM SEA EL LSB DE LA CUENTA 
	              CUENTA(1) WHEN "01", --ELEGIMOS QUE LA SALIDA DEL PWM SEA EL BIT 1 DE LA CUENTA 
					  CUENTA(2) WHEN "10", --ELEGIMOS QUE LA SALIDA DEL PWM SEA EL BIT 2 DE LA CUENTA
					  CUENTA(3) WHEN OTHERS; --ELEGIMOS QUE LA SALIDA DEL PWM SEA EL MSB DE LA CUENTA 
END MODULACION;