LIBRARY IEEE; 

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 

ENTITY POR_DOS IS 
PORT
(
	ENTRADA1, ENTRADA2 : IN BIT;
	SELECTOR : IN STD_LOGIC_VECTOR(1 DOWNTO 0); --En este caso el selector tiene 2 bits para poder elegir mas opciones 
	SALIDA1: OUT BIT
);
END POR_DOS;

ARCHITECTURE SELECTOR_DOBLE OF POR_DOS IS 
BEGIN 
WITH SELECTOR SELECT 
SALIDA1 <= ENTRADA1 OR ENTRADA2 WHEN "00",
          ENTRADA1 AND ENTRADA2 WHEN "01",
			 ENTRADA1 XOR ENTRADA2 WHEN "10",
			 ENTRADA2 XNOR ENTRADA1	 WHEN OTHERS;
END SELECTOR_DOBLE;